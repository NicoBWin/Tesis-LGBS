
// 48M clk
`define BAUD8M_CLK48M 6
`define BAUD8M_CLK48M 2

// 24M clk
`define BAUD8M_CLK24M 3
`define BAUD24M_CLK24M 1