// 48M clk
`define BAUD6M_CLK48M 4'd4
`define BAUD1M_CLK48M 5'd24

// 24M clk
`define BAUD1M_CLK24M 4'd12
`define BAUD4M_CLK24M 4'd3
`define BAUD6M_CLK24M 4'd2
`define BAUD12M_CLK24M 4'd1

// 12M clk
`define BAUD6M_CLK12M 4'd1
