
// 48Mhz
`define RATE4M8_CLK48M 10