
// 24M clk

`define BAUD8M 3
`define BAUD24M 1