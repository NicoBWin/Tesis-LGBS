// 48M clk
`define BAUD6M_CLK48M 4'd4
`define BAUD3M_CLK48M 4'd8
`define BAUD1M_CLK48M 5'd24
`define BAUD115200_CLK48M 10'd417

// 24M clk
`define BAUD1M_CLK24M 4'd12
`define BAUD4M_CLK24M 4'd3
`define BAUD6M_CLK24M 4'd2
`define BAUD12M_CLK24M 4'd1

// 12M clk
`define BAUD6M_CLK12M 4'd1
