
// 24Mhz
`define SAMPLE240K_CLK24M 100