
// 48Mhz
`define RATE2M4_CLK48M 10
`define RATE4M8_CLK48M 5

// 24Mhz
`define RATE250k_CLK24M 48
`define RATE1M2_CLK24M 10
`define RATE2M4_CLK24M 5
`define RATE3M_CLK24M 4
`define RATE4M_CLK24M 3
`define RATE6M_CLK24M 2
`define RATE12M_CLK24M 1
