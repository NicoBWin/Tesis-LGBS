
module generator();

    

endmodule