
// 24Mhz
`define MSEC_10 240000
`define MSEC_100 2400000
`define MSEC_500 12000000
`define SEC_1 24000000  // Contador de 1 segundo con un reloj de 48Mhz
`define SEC_2 48000000  // Contador de 2 segundos con un reloj de 48Mhz
`define SEC_5 120000000 // Contador de 5 segundos con un reloj de 48Mhz