
`define SAMPLE1M2 20