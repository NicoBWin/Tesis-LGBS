/*
    Este module se encarga de generar las señales de SPWM que se enviaran 
    a cada uno de los submodulos FPGA_modulo. Tambien enviara la señal de disparo para
    sincronizarlos.  
*/

module top(
    input wire gpio_25,

    output wire led_green,
    output wire led_red,
    output wire led_blue,
    output wire gpio_23,
    output wire gpio_26,
    output wire gpio_27,
    output wire gpio_32,
);

/*
*******************
*   Ports setup   *
*******************
*/

    wire tx;
    wire rx;
    wire tx_busy;
    wire rx_done;
    wire parity_error;
    
    assign tx = gpio_23;
    assign rx = gpio_25;
    assign tx_busy = gpio_26;
    assign rx_done = gpio_27;
    assign parity_error = gpio_32;
/*
*********************
*   HFClock setup   *
*********************
*/  
    wire clk;
    SB_HFOSC  #(.CLKHF_DIV("0b11") // 48 MHz = ~48 MHz / 1 (0b00=1, 0b01=2, 0b10=4, 0b11=8)
    )  
    hf_osc (.CLKHFPU(1'b1), .CLKHFEN(1'b1), .CLKHF(clk));

/*
*****************************
*   Variables declaration   *
*****************************
*/  
    localparam turn_on = 8'b10101010;
    localparam turn_off = 8'b01010101;
    localparam toggle = 8'b11000011;
    localparam OFF = 1;
    localparam ON = 0;

    wire [7:0] data_received;
    wire start_tx;

    reg [7:0] data_to_tx = toggle;
    reg reset = 0;
/*
*************************************
*   External Modules declarations   *
*************************************
*/

    uart_tx transmitter(
        .clk(clk), 
        .reset(reset), 
        .data_to_tx(data_to_tx), 
        .start_tx(start_tx), 
        .tx(tx), 
        .tx_busy(tx_busy)
    );

    uart_rx receiver(
        .clk(clk), 
        .reset(reset), 
        .rx(rx),
        .data_received(data_received), 
        .rx_done(rx_done), 
        .parity_error(parity_error)
    );

/*
******************
*   Statements   *
******************
*/

    parameter INIT  = 3'b001; 
    parameter UART_SEND = 3'b010; 
    parameter END_TX = 3'b100;
    parameter WAIT = 3'b101;

    reg led_r = OFF;
    reg led_g = OFF;
    reg led_b = OFF;
    reg[2:0] state = INIT;
    reg[31:0] counter = 0;

    assign led_red = led_r;
    assign led_green = led_g;
    assign led_blue = led_b;

    always @(posedge clk) begin
        case (state)

            INIT: begin
                reset   <= 1;
                led_r   <= OFF;
                led_g   <= OFF;
                led_b   <= OFF;
                counter <= counter + 1;
                if (counter >= 6000000) begin
                    reset <= 0;
                    state <= UART_SEND;
                    counter <= 0;
                end
            end

            UART_SEND: begin
                led_b   <= ON;
                start_tx <= 1;

                if (rx_done)
                    if (data_received == data_to_tx) begin
                        led_r <= ~led_r;
                        counter <= 0;
                    end
                    else begin
                        led_r <= OFF;
                    end
                else
                    counter <= counter + 1;

                if (counter >= 10*6000000) begin
                    start_tx <= 0;
                    state <= END_TX;
                    counter <= 0;
                end
            end

            END_TX: begin
                led_b <= OFF;         // Turn off green LED
                state <= WAIT;        // Move to waiting state
                counter <= 0;
            end

            WAIT: begin
                counter <= counter + 1;
                if (counter >= 6000000) begin
                    state <= INIT;    // Restart the cycle
                    counter <= 0;
                end
            end

        endcase
    end

endmodule