
// 48M clk
`define BAUD8M 6
`define BAUD24M 2