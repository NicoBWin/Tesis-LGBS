
`define UP 0
`define DOWN 1
`define FREC240K 10
