
// 48Mhz
`define MSEC_10 480000
`define MSEC_100 4800000
`define MSEC_500 24000000
`define SEC_1 48000000  // Contador de 1 segundo con un reloj de 48Mhz
`define SEC_2 96000000  // Contador de 2 segundos con un reloj de 48Mhz
`define SEC_5 240000000 // Contador de 5 segundos con un reloj de 48Mhz