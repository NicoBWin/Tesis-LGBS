// 24M clk
`define BAUD1M_CLK24M 12
`define BAUD4M_CLK24M 3
`define BAUD6M_CLK24M 2
`define BAUD12M_CLK24M 1

// 12M clk
`define BAUD6M_CLK12M 1
