
// SPI codes
`define PIPE_MODE 16'hB0CA